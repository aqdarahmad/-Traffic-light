module cla(sum,cout,a,b,cin);
output [5:0]sum;output cout;
input [5:0]a,b; input cin;
wire p0,p1,p2,p3,p4,p5,g0,g1,g2,g3,g4,g5,c1,c2,c3,c4,c5,c6 ;
wire w1,w2,w3,w4,w5,w6,w7,w8,w9,w10;
wire c44,e1,e2,e3,e4,e5,e11,e22,e33,e44,e55,e9;
xor #10 (p0,a[0],b[0]); xor #10 (p1,a[1],b[1]);
xor #10(p2,a[2],b[2]);xor #10(p3,a[3],b[3]);
xor #10(p4,a[4],b[4]); xor #10(p5,a[5],b[5]);
and #10 (g0,a[0],b[0]);and #10 (g1,a[1],b[1]);
and #10 (g2,a[2],b[2]); and #10 (g3,a[3],b[3]);
and #10 (g4,a[4],b[4]); and #10 (g5,a[5],b[5]);
assign c0=cin;
and #10(w1,p0,cin); or #10(c1,w1,g0);and #10(w2,p1,g0);
and #10(w3,p1,p0,cin); or #10(c2,w3,w2,g1);
and #10 (w4,p2,g1);and #10(w5,p2,p1,g0);
and #10(w6,p1,p0,cin); or#10(c3,w6,w5,w4,g2);
and #10(w7,p3,g2);and #10(w8,p3,p2,g1);and #10 (w9,p3,p2,p1,g0);
and #10 (w10,p3,p2,p1,p0,cin); or #10(c4,w10,w9,w8,w7,cin);
and #10(e1,p4,g3);and #10 (e2,p4,p3,g2);
and #10 (e3,p4,p3,p2,g1);and #10 (e4,p4,p3,p2,p1,p0,cin);
and #10 (e5,p4,p3,p2,p1,g0);or #10 (c5,g4,e1,e2,e3,e4,e5);
and #10(e11,p5,g4);and #10 (e22,p5,p4,p3,g2);
and #10 (e9,p5,p4,p3,p2,g1);and #10 (e33,p5,p4,g3);
and #10 (e44,p5,p4,p3,p2,p1,p0,cin);
and #10 (e55,p5,p4,p3,p2,p1,g0);
or #10 (c6,g5,e11,e22,e9,e33,e44,e55);xor #10(sum[0],p0,c0);
xor #10(sum[1],p1,c1); xor #10(sum[2],p2,c2);
xor #10(sum[3],p3,c3);xor #10(sum[4],p4,c5);
xor #10(sum[5],p5,c6);assign cout=c4;
endmodule
